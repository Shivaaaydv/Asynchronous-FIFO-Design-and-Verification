// File: /master/fifo_wsqr.sv
// Description: Defines the sequencer typedef for asynchronous fifo transactions.
// Author: Karankumar Nevage | Email: karanpr9423@gmail.com
// Version: 0.1
//==================================================================================================================================================
typedef uvm_sequencer#(fifo_tx) fifo_wsqr;
//==================================================================================================================================================
