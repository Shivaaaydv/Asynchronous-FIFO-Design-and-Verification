// File: /master/fifo_rsqr.sv
// Description: Defines the read sequencer typedef for asynchronous fifo transactions.
// Author: Karankumar Nevage | Email: karanpr9423@gmail.com
// Version: 0.1
//==================================================================================================================================================
typedef uvm_sequencer#(fifo_tx) fifo_rsqr;
//==================================================================================================================================================
